11111111111
22222222222
add 3333333
add 2222222
