11111111111
add 2222222
